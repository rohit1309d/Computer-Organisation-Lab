$date
   Thu Sep 17 23:38:08 2020
$end
$version
  2020.1
$end
$timescale
  1ps
$end
$scope module serial_adder_tb $end
$var reg 4 ! data_a [3:0] $end
$var reg 4 " data_b [3:0] $end
$var reg 1 # clk $end
$var wire 4 $ sum [3:0] $end
$var wire 1 % cout $end
$scope module s_adder $end
$var wire 4 & data_a [3:0] $end
$var wire 4 ' data_b [3:0] $end
$var wire 1 ( clk $end
$var reg 4 ) sum [3:0] $end
$var reg 3 * count [2:0] $end
$var reg 1 + cout $end
$var wire 1 , wire_a $end
$var wire 1 - wire_b $end
$var wire 1 . cout_temp $end
$var wire 1 / cin $end
$var wire 1 0 s $end
$scope module piso_a $end
$var wire 1 ( clk $end
$var wire 4 & data [3:0] $end
$var reg 1 1 out $end
$var reg 4 2 memory [3:0] $end
$upscope $end
$scope module piso_b $end
$var wire 1 ( clk $end
$var wire 4 ' data [3:0] $end
$var reg 1 3 out $end
$var reg 4 4 memory [3:0] $end
$upscope $end
$scope module adder $end
$var wire 1 , a $end
$var wire 1 - b $end
$var wire 1 / cin $end
$var wire 1 0 sum $end
$var wire 1 . cout $end
$upscope $end
$scope module dff $end
$var wire 1 . d $end
$var wire 1 ( clk $end
$var reg 1 5 out $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
b10 !
b10 "
0#
bx $
x%
b10 &
b10 '
0(
bx )
bx *
x+
x,
x-
x.
x/
x0
x1
bx 2
x3
bx 4
x5
$end
#10000
1#
bx $
1(
bx )
x+
x1
b0xxx 2
x3
b0xxx 4
x5
#20000
0#
0(
#30000
1#
bx $
1(
bx )
x+
x1
b0xx 2
x3
b0xx 4
x5
#40000
0#
0(
#50000
1#
bx $
1(
bx )
x+
x1
b0x 2
x3
b0x 4
x5
#60000
0#
0(
#70000
1#
bx $
1(
bx )
x+
x1
b0 2
x3
b0 4
x5
#80000
0#
0(
#90000
1#
bx $
1(
bx )
x+
0,
0-
0.
01
03
x5
#100000
0#
0(
#110000
1#
bx $
0%
1(
bx )
0+
0/
00
01
03
05
#120000
0#
0(
#130000
1#
b0xxx $
1(
b0xxx )
0+
01
03
05
#140000
0#
0(
#150000
1#
b0xx $
1(
b0xx )
0+
01
03
05
#160000
0#
0(
#170000
1#
b0x $
1(
b0x )
0+
01
03
05
#180000
0#
0(
#190000
1#
b0 $
1(
b0 )
0+
01
03
05
#200000
b100 !
b101 "
0#
b100 &
b101 '
0(
#210000
1#
1(
b0 )
0+
01
03
05
#220000
0#
0(
#230000
1#
1(
b0 )
0+
01
03
05
#240000
0#
0(
#250000
1#
1(
b0 )
0+
01
03
05
#260000
0#
0(
#270000
1#
1(
b0 )
0+
01
03
05
#280000
0#
0(
#290000
1#
1(
b0 )
0+
01
03
05
#300000
0#
0(
#310000
1#
1(
b0 )
0+
01
03
05
#320000
0#
0(
#330000
1#
1(
b0 )
0+
01
03
05
#340000
0#
0(
#350000
1#
1(
b0 )
0+
01
03
05
#360000
0#
0(
#370000
1#
1(
b0 )
0+
01
03
05
#380000
0#
0(
#390000
1#
1(
b0 )
0+
01
03
05
